library verilog;
use verilog.vl_types.all;
entity JK_async_sync_tb is
end JK_async_sync_tb;

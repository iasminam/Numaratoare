library verilog;
use verilog.vl_types.all;
entity JK_sync_counter_tb is
end JK_sync_counter_tb;

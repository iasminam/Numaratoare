library verilog;
use verilog.vl_types.all;
entity JK_async_counter_tb is
end JK_async_counter_tb;
